VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mpw2304c_mp
  CLASS BLOCK ;
  FOREIGN mpw2304c_mp ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.005 BY 0.005 ;
END mpw2304c_mp
END LIBRARY

